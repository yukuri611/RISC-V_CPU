`ifndef DEFINES_VH
`define DEFINES_VH

`define OP_OP_IMM 7'b0010011
`define OP_OP     7'b0110011

`endif
