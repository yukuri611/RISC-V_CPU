`ifndef DEFINES_VH
`define DEFINES_VH

`define OP_IMM    7'b0010011
`define OP_LOAD   7'b0000011
`define OP_STORE  7'b0100011
`define OP_R_TYPE 7'b0110011
`define OP_BRANCH 7'b1100011
`endif
