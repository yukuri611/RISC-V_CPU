`ifndef DEFINES_VH
`define DEFINES_VH

`define OP_IMM    7'b0010011
`define OP_LOAD   7'b0000011
`define OP_STORE  7'b0100011

`endif
